----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    14:12:55 02/06/2024 
-- Design Name: 
-- Module Name:    moi_top_modul - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity top_modul is
port(
	clk: in std_logic;
	led: out std_logic_vector(7 downto 0);
	switch: in std_logic_vector(2 downto 0);
	--SPI DAC
	nSync : out std_logic;
	CLK_DAC : out std_logic;
	D1  : out std_logic;
	D2  : out std_logic;
	--ADC
	nSync_ADC : out std_logic;
	CLK_ADC : out std_logic;
	DataADC : in std_logic;
	DataADC2 : in std_logic
);
end top_modul;

architecture Behavioral of top_modul is

signal cnt: integer range 0 to 1151:=0;--make it a constant
signal clk_da2: std_logic;
signal pila: integer range 0 to 4095:=0;
signal ink: integer range 0 to 1:=1;
signal ADC: std_logic_vector(11 downto 0);
signal ADC1: std_logic_vector(11 downto 0);
signal RES_out: std_logic_vector(11 downto 0);
signal Data1: std_logic_vector(11 DOWNTO 0);
signal Data2: std_logic_vector(11 DOWNTO 0);
signal i: integer range 0 to 4095:=0;
type ROM_array is array(0 to 4095)of integer;
constant sin_array: ROM_array:= (
0 => 2048,
1 => 2113,
2 => 2179,
3 => 2245,
4 => 2311,
5 => 2377,
6 => 2443,
7 => 2509,
8 => 2575,
9 => 2641,
10 => 2707,
11 => 2773,
12 => 2839,
13 => 2905,
14 => 2971,
15 => 3037,
16 => 3103,
17 => 3169,
18 => 3235,
19 => 3301,
20 => 3366,
21 => 3432,
22 => 3498,
23 => 3564,
24 => 3630,
25 => 3696,
26 => 3762,
27 => 3828,
28 => 3894,
29 => 3960,
30 => 4026,
31 => 4091,
32 => 4157,
33 => 4223,
34 => 4289,
35 => 4355,
36 => 4421,
37 => 4487,
38 => 4552,
39 => 4618,
40 => 4684,
41 => 4750,
42 => 4816,
43 => 4882,
44 => 4947,
45 => 5013,
46 => 5079,
47 => 5145,
48 => 5211,
49 => 5276,
50 => 5342,
51 => 5408,
52 => 5474,
53 => 5539,
54 => 5605,
55 => 5671,
56 => 5737,
57 => 5802,
58 => 5868,
59 => 5934,
60 => 5999,
61 => 6065,
62 => 6131,
63 => 6196,
64 => 6262,
65 => 6328,
66 => 6393,
67 => 6459,
68 => 6524,
69 => 6590,
70 => 6656,
71 => 6721,
72 => 6787,
73 => 6852,
74 => 6918,
75 => 6983,
76 => 7049,
77 => 7114,
78 => 7180,
79 => 7245,
80 => 7311,
81 => 7376,
82 => 7442,
83 => 7507,
84 => 7573,
85 => 7638,
86 => 7703,
87 => 7769,
88 => 7834,
89 => 7899,
90 => 7965,
91 => 8030,
92 => 8095,
93 => 8161,
94 => 8226,
95 => 8291,
96 => 8357,
97 => 8422,
98 => 8487,
99 => 8552,
100 => 8617,
101 => 8683,
102 => 8748,
103 => 8813,
104 => 8878,
105 => 8943,
106 => 9008,
107 => 9073,
108 => 9138,
109 => 9203,
110 => 9268,
111 => 9333,
112 => 9398,
113 => 9463,
114 => 9528,
115 => 9593,
116 => 9658,
117 => 9723,
118 => 9788,
119 => 9853,
120 => 9918,
121 => 9983,
122 => 10047,
123 => 10112,
124 => 10177,
125 => 10242,
126 => 10306,
127 => 10371,
128 => 10436,
129 => 10501,
130 => 10565,
131 => 10630,
132 => 10694,
133 => 10759,
134 => 10824,
135 => 10888,
136 => 10953,
137 => 11017,
138 => 11082,
139 => 11146,
140 => 11211,
141 => 11275,
142 => 11340,
143 => 11404,
144 => 11468,
145 => 11533,
146 => 11597,
147 => 11661,
148 => 11726,
149 => 11790,
150 => 11854,
151 => 11918,
152 => 11982,
153 => 12047,
154 => 12111,
155 => 12175,
156 => 12239,
157 => 12303,
158 => 12367,
159 => 12431,
160 => 12495,
161 => 12559,
162 => 12623,
163 => 12687,
164 => 12751,
165 => 12815,
166 => 12878,
167 => 12942,
168 => 13006,
169 => 13070,
170 => 13134,
171 => 13197,
172 => 13261,
173 => 13325,
174 => 13388,
175 => 13452,
176 => 13515,
177 => 13579,
178 => 13643,
179 => 13706,
180 => 13770,
181 => 13833,
182 => 13896,
183 => 13960,
184 => 14023,
185 => 14086,
186 => 14150,
187 => 14213,
188 => 14276,
189 => 14340,
190 => 14403,
191 => 14466,
192 => 14529,
193 => 14592,
194 => 14655,
195 => 14718,
196 => 14781,
197 => 14844,
198 => 14907,
199 => 14970,
200 => 15033,
201 => 15096,
202 => 15159,
203 => 15221,
204 => 15284,
205 => 15347,
206 => 15410,
207 => 15472,
208 => 15535,
209 => 15598,
210 => 15660,
211 => 15723,
212 => 15785,
213 => 15848,
214 => 15910,
215 => 15973,
216 => 16035,
217 => 16097,
218 => 16160,
219 => 16222,
220 => 16284,
221 => 16346,
222 => 16409,
223 => 16471,
224 => 16533,
225 => 16595,
226 => 16657,
227 => 16719,
228 => 16781,
229 => 16843,
230 => 16905,
231 => 16967,
232 => 17029,
233 => 17090,
234 => 17152,
235 => 17214,
236 => 17276,
237 => 17337,
238 => 17399,
239 => 17461,
240 => 17522,
241 => 17584,
242 => 17645,
243 => 17707,
244 => 17768,
245 => 17829,
246 => 17891,
247 => 17952,
248 => 18013,
249 => 18074,
250 => 18136,
251 => 18197,
252 => 18258,
253 => 18319,
254 => 18380,
255 => 18441,
256 => 18502,
257 => 18563,
258 => 18624,
259 => 18685,
260 => 18745,
261 => 18806,
262 => 18867,
263 => 18928,
264 => 18988,
265 => 19049,
266 => 19109,
267 => 19170,
268 => 19230,
269 => 19291,
270 => 19351,
271 => 19412,
272 => 19472,
273 => 19532,
274 => 19592,
275 => 19653,
276 => 19713,
277 => 19773,
278 => 19833,
279 => 19893,
280 => 19953,
281 => 20013,
282 => 20073,
283 => 20133,
284 => 20192,
285 => 20252,
286 => 20312,
287 => 20372,
288 => 20431,
289 => 20491,
290 => 20550,
291 => 20610,
292 => 20669,
293 => 20729,
294 => 20788,
295 => 20848,
296 => 20907,
297 => 20966,
298 => 21025,
299 => 21085,
300 => 21144,
301 => 21203,
302 => 21262,
303 => 21321,
304 => 21380,
305 => 21439,
306 => 21497,
307 => 21556,
308 => 21615,
309 => 21674,
310 => 21732,
311 => 21791,
312 => 21850,
313 => 21908,
314 => 21967,
315 => 22025,
316 => 22083,
317 => 22142,
318 => 22200,
319 => 22258,
320 => 22316,
321 => 22375,
322 => 22433,
323 => 22491,
324 => 22549,
325 => 22607,
326 => 22665,
327 => 22722,
328 => 22780,
329 => 22838,
330 => 22896,
331 => 22953,
332 => 23011,
333 => 23069,
334 => 23126,
335 => 23183,
336 => 23241,
337 => 23298,
338 => 23356,
339 => 23413,
340 => 23470,
341 => 23527,
342 => 23584,
343 => 23641,
344 => 23698,
345 => 23755,
346 => 23812,
347 => 23869,
348 => 23926,
349 => 23983,
350 => 24039,
351 => 24096,
352 => 24153,
353 => 24209,
354 => 24266,
355 => 24322,
356 => 24379,
357 => 24435,
358 => 24491,
359 => 24547,
360 => 24604,
361 => 24660,
362 => 24716,
363 => 24772,
364 => 24828,
365 => 24884,
366 => 24940,
367 => 24995,
368 => 25051,
369 => 25107,
370 => 25162,
371 => 25218,
372 => 25274,
373 => 25329,
374 => 25384,
375 => 25440,
376 => 25495,
377 => 25550,
378 => 25606,
379 => 25661,
380 => 25716,
381 => 25771,
382 => 25826,
383 => 25881,
384 => 25936,
385 => 25990,
386 => 26045,
387 => 26100,
388 => 26155,
389 => 26209,
390 => 26264,
391 => 26318,
392 => 26373,
393 => 26427,
394 => 26481,
395 => 26535,
396 => 26590,
397 => 26644,
398 => 26698,
399 => 26752,
400 => 26806,
401 => 26860,
402 => 26914,
403 => 26967,
404 => 27021,
405 => 27075,
406 => 27128,
407 => 27182,
408 => 27235,
409 => 27289,
410 => 27342,
411 => 27395,
412 => 27449,
413 => 27502,
414 => 27555,
415 => 27608,
416 => 27661,
417 => 27714,
418 => 27767,
419 => 27820,
420 => 27873,
421 => 27925,
422 => 27978,
423 => 28030,
424 => 28083,
425 => 28135,
426 => 28188,
427 => 28240,
428 => 28292,
429 => 28345,
430 => 28397,
431 => 28449,
432 => 28501,
433 => 28553,
434 => 28605,
435 => 28657,
436 => 28708,
437 => 28760,
438 => 28812,
439 => 28863,
440 => 28915,
441 => 28966,
442 => 29018,
443 => 29069,
444 => 29120,
445 => 29172,
446 => 29223,
447 => 29274,
448 => 29325,
449 => 29376,
450 => 29427,
451 => 29477,
452 => 29528,
453 => 29579,
454 => 29630,
455 => 29680,
456 => 29731,
457 => 29781,
458 => 29831,
459 => 29882,
460 => 29932,
461 => 29982,
462 => 30032,
463 => 30082,
464 => 30132,
465 => 30182,
466 => 30232,
467 => 30282,
468 => 30332,
469 => 30381,
470 => 30431,
471 => 30480,
472 => 30530,
473 => 30579,
474 => 30628,
475 => 30678,
476 => 30727,
477 => 30776,
478 => 30825,
479 => 30874,
480 => 30923,
481 => 30972,
482 => 31020,
483 => 31069,
484 => 31118,
485 => 31166,
486 => 31215,
487 => 31263,
488 => 31312,
489 => 31360,
490 => 31408,
491 => 31456,
492 => 31504,
493 => 31552,
494 => 31600,
495 => 31648,
496 => 31696,
497 => 31744,
498 => 31791,
499 => 31839,
500 => 31887,
501 => 31934,
502 => 31981,
503 => 32029,
504 => 32076,
505 => 32123,
506 => 32170,
507 => 32217,
508 => 32264,
509 => 32311,
510 => 32358,
511 => 32405,
512 => 32451,
513 => 32498,
514 => 32544,
515 => 32591,
516 => 32637,
517 => 32684,
518 => 32730,
519 => 32776,
520 => 32822,
521 => 32868,
522 => 32914,
523 => 32960,
524 => 33006,
525 => 33052,
526 => 33097,
527 => 33143,
528 => 33188,
529 => 33234,
530 => 33279,
531 => 33324,
532 => 33370,
533 => 33415,
534 => 33460,
535 => 33505,
536 => 33550,
537 => 33595,
538 => 33639,
539 => 33684,
540 => 33729,
541 => 33773,
542 => 33818,
543 => 33862,
544 => 33907,
545 => 33951,
546 => 33995,
547 => 34039,
548 => 34083,
549 => 34127,
550 => 34171,
551 => 34215,
552 => 34258,
553 => 34302,
554 => 34346,
555 => 34389,
556 => 34433,
557 => 34476,
558 => 34519,
559 => 34562,
560 => 34606,
561 => 34649,
562 => 34692,
563 => 34734,
564 => 34777,
565 => 34820,
566 => 34863,
567 => 34905,
568 => 34948,
569 => 34990,
570 => 35033,
571 => 35075,
572 => 35117,
573 => 35159,
574 => 35201,
575 => 35243,
576 => 35285,
577 => 35327,
578 => 35369,
579 => 35410,
580 => 35452,
581 => 35493,
582 => 35535,
583 => 35576,
584 => 35617,
585 => 35658,
586 => 35700,
587 => 35741,
588 => 35781,
589 => 35822,
590 => 35863,
591 => 35904,
592 => 35944,
593 => 35985,
594 => 36025,
595 => 36066,
596 => 36106,
597 => 36146,
598 => 36186,
599 => 36227,
600 => 36266,
601 => 36306,
602 => 36346,
603 => 36386,
604 => 36426,
605 => 36465,
606 => 36505,
607 => 36544,
608 => 36583,
609 => 36623,
610 => 36662,
611 => 36701,
612 => 36740,
613 => 36779,
614 => 36818,
615 => 36856,
616 => 36895,
617 => 36934,
618 => 36972,
619 => 37011,
620 => 37049,
621 => 37087,
622 => 37125,
623 => 37164,
624 => 37202,
625 => 37240,
626 => 37277,
627 => 37315,
628 => 37353,
629 => 37390,
630 => 37428,
631 => 37465,
632 => 37503,
633 => 37540,
634 => 37577,
635 => 37614,
636 => 37651,
637 => 37688,
638 => 37725,
639 => 37762,
640 => 37799,
641 => 37835,
642 => 37872,
643 => 37908,
644 => 37945,
645 => 37981,
646 => 38017,
647 => 38053,
648 => 38089,
649 => 38125,
650 => 38161,
651 => 38197,
652 => 38232,
653 => 38268,
654 => 38303,
655 => 38339,
656 => 38374,
657 => 38409,
658 => 38444,
659 => 38480,
660 => 38515,
661 => 38549,
662 => 38584,
663 => 38619,
664 => 38654,
665 => 38688,
666 => 38723,
667 => 38757,
668 => 38791,
669 => 38826,
670 => 38860,
671 => 38894,
672 => 38928,
673 => 38962,
674 => 38995,
675 => 39029,
676 => 39063,
677 => 39096,
678 => 39130,
679 => 39163,
680 => 39196,
681 => 39229,
682 => 39262,
683 => 39295,
684 => 39328,
685 => 39361,
686 => 39394,
687 => 39427,
688 => 39459,
689 => 39492,
690 => 39524,
691 => 39556,
692 => 39588,
693 => 39621,
694 => 39653,
695 => 39684,
696 => 39716,
697 => 39748,
698 => 39780,
699 => 39811,
700 => 39843,
701 => 39874,
702 => 39906,
703 => 39937,
704 => 39968,
705 => 39999,
706 => 40030,
707 => 40061,
708 => 40092,
709 => 40122,
710 => 40153,
711 => 40183,
712 => 40214,
713 => 40244,
714 => 40274,
715 => 40305,
716 => 40335,
717 => 40365,
718 => 40394,
719 => 40424,
720 => 40454,
721 => 40484,
722 => 40513,
723 => 40542,
724 => 40572,
725 => 40601,
726 => 40630,
727 => 40659,
728 => 40688,
729 => 40717,
730 => 40746,
731 => 40775,
732 => 40803,
733 => 40832,
734 => 40860,
735 => 40889,
736 => 40917,
737 => 40945,
738 => 40973,
739 => 41001,
740 => 41029,
741 => 41057,
742 => 41084,
743 => 41112,
744 => 41139,
745 => 41167,
746 => 41194,
747 => 41221,
748 => 41249,
749 => 41276,
750 => 41303,
751 => 41329,
752 => 41356,
753 => 41383,
754 => 41410,
755 => 41436,
756 => 41462,
757 => 41489,
758 => 41515,
759 => 41541,
760 => 41567,
761 => 41593,
762 => 41619,
763 => 41645,
764 => 41670,
765 => 41696,
766 => 41721,
767 => 41747,
768 => 41772,
769 => 41797,
770 => 41822,
771 => 41847,
772 => 41872,
773 => 41897,
774 => 41922,
775 => 41946,
776 => 41971,
777 => 41995,
778 => 42020,
779 => 42044,
780 => 42068,
781 => 42092,
782 => 42116,
783 => 42140,
784 => 42164,
785 => 42188,
786 => 42211,
787 => 42235,
788 => 42258,
789 => 42281,
790 => 42305,
791 => 42328,
792 => 42351,
793 => 42374,
794 => 42397,
795 => 42419,
796 => 42442,
797 => 42464,
798 => 42487,
799 => 42509,
800 => 42532,
801 => 42554,
802 => 42576,
803 => 42598,
804 => 42620,
805 => 42641,
806 => 42663,
807 => 42685,
808 => 42706,
809 => 42728,
810 => 42749,
811 => 42770,
812 => 42791,
813 => 42812,
814 => 42833,
815 => 42854,
816 => 42875,
817 => 42895,
818 => 42916,
819 => 42936,
820 => 42957,
821 => 42977,
822 => 42997,
823 => 43017,
824 => 43037,
825 => 43057,
826 => 43077,
827 => 43097,
828 => 43116,
829 => 43136,
830 => 43155,
831 => 43174,
832 => 43194,
833 => 43213,
834 => 43232,
835 => 43251,
836 => 43269,
837 => 43288,
838 => 43307,
839 => 43325,
840 => 43344,
841 => 43362,
842 => 43380,
843 => 43398,
844 => 43416,
845 => 43434,
846 => 43452,
847 => 43470,
848 => 43487,
849 => 43505,
850 => 43522,
851 => 43540,
852 => 43557,
853 => 43574,
854 => 43591,
855 => 43608,
856 => 43625,
857 => 43642,
858 => 43658,
859 => 43675,
860 => 43692,
861 => 43708,
862 => 43724,
863 => 43740,
864 => 43756,
865 => 43772,
866 => 43788,
867 => 43804,
868 => 43820,
869 => 43835,
870 => 43851,
871 => 43866,
872 => 43881,
873 => 43897,
874 => 43912,
875 => 43927,
876 => 43942,
877 => 43956,
878 => 43971,
879 => 43986,
880 => 44000,
881 => 44015,
882 => 44029,
883 => 44043,
884 => 44057,
885 => 44071,
886 => 44085,
887 => 44099,
888 => 44113,
889 => 44126,
890 => 44140,
891 => 44153,
892 => 44167,
893 => 44180,
894 => 44193,
895 => 44206,
896 => 44219,
897 => 44232,
898 => 44244,
899 => 44257,
900 => 44269,
901 => 44282,
902 => 44294,
903 => 44306,
904 => 44319,
905 => 44331,
906 => 44343,
907 => 44354,
908 => 44366,
909 => 44378,
910 => 44389,
911 => 44401,
912 => 44412,
913 => 44423,
914 => 44434,
915 => 44445,
916 => 44456,
917 => 44467,
918 => 44478,
919 => 44488,
920 => 44499,
921 => 44509,
922 => 44520,
923 => 44530,
924 => 44540,
925 => 44550,
926 => 44560,
927 => 44570,
928 => 44580,
929 => 44589,
930 => 44599,
931 => 44608,
932 => 44618,
933 => 44627,
934 => 44636,
935 => 44645,
936 => 44654,
937 => 44663,
938 => 44671,
939 => 44680,
940 => 44689,
941 => 44697,
942 => 44705,
943 => 44714,
944 => 44722,
945 => 44730,
946 => 44738,
947 => 44745,
948 => 44753,
949 => 44761,
950 => 44768,
951 => 44776,
952 => 44783,
953 => 44790,
954 => 44797,
955 => 44804,
956 => 44811,
957 => 44818,
958 => 44825,
959 => 44831,
960 => 44838,
961 => 44844,
962 => 44851,
963 => 44857,
964 => 44863,
965 => 44869,
966 => 44875,
967 => 44881,
968 => 44886,
969 => 44892,
970 => 44898,
971 => 44903,
972 => 44908,
973 => 44913,
974 => 44919,
975 => 44924,
976 => 44928,
977 => 44933,
978 => 44938,
979 => 44943,
980 => 44947,
981 => 44951,
982 => 44956,
983 => 44960,
984 => 44964,
985 => 44968,
986 => 44972,
987 => 44976,
988 => 44979,
989 => 44983,
990 => 44987,
991 => 44990,
992 => 44993,
993 => 44996,
994 => 44999,
995 => 45002,
996 => 45005,
997 => 45008,
998 => 45011,
999 => 45013,
1000 => 45016,
1001 => 45018,
1002 => 45021,
1003 => 45023,
1004 => 45025,
1005 => 45027,
1006 => 45029,
1007 => 45030,
1008 => 45032,
1009 => 45034,
1010 => 45035,
1011 => 45036,
1012 => 45038,
1013 => 45039,
1014 => 45040,
1015 => 45041,
1016 => 45042,
1017 => 45043,
1018 => 45043,
1019 => 45044,
1020 => 45044,
1021 => 45045,
1022 => 45045,
1023 => 45045,
1024 => 45045,
1025 => 45045,
1026 => 45045,
1027 => 45045,
1028 => 45044,
1029 => 45044,
1030 => 45043,
1031 => 45043,
1032 => 45042,
1033 => 45041,
1034 => 45040,
1035 => 45039,
1036 => 45038,
1037 => 45036,
1038 => 45035,
1039 => 45034,
1040 => 45032,
1041 => 45030,
1042 => 45029,
1043 => 45027,
1044 => 45025,
1045 => 45023,
1046 => 45021,
1047 => 45018,
1048 => 45016,
1049 => 45013,
1050 => 45011,
1051 => 45008,
1052 => 45005,
1053 => 45002,
1054 => 44999,
1055 => 44996,
1056 => 44993,
1057 => 44990,
1058 => 44987,
1059 => 44983,
1060 => 44979,
1061 => 44976,
1062 => 44972,
1063 => 44968,
1064 => 44964,
1065 => 44960,
1066 => 44956,
1067 => 44951,
1068 => 44947,
1069 => 44943,
1070 => 44938,
1071 => 44933,
1072 => 44928,
1073 => 44924,
1074 => 44919,
1075 => 44913,
1076 => 44908,
1077 => 44903,
1078 => 44898,
1079 => 44892,
1080 => 44886,
1081 => 44881,
1082 => 44875,
1083 => 44869,
1084 => 44863,
1085 => 44857,
1086 => 44851,
1087 => 44844,
1088 => 44838,
1089 => 44831,
1090 => 44825,
1091 => 44818,
1092 => 44811,
1093 => 44804,
1094 => 44797,
1095 => 44790,
1096 => 44783,
1097 => 44776,
1098 => 44768,
1099 => 44761,
1100 => 44753,
1101 => 44745,
1102 => 44738,
1103 => 44730,
1104 => 44722,
1105 => 44714,
1106 => 44705,
1107 => 44697,
1108 => 44689,
1109 => 44680,
1110 => 44671,
1111 => 44663,
1112 => 44654,
1113 => 44645,
1114 => 44636,
1115 => 44627,
1116 => 44618,
1117 => 44608,
1118 => 44599,
1119 => 44589,
1120 => 44580,
1121 => 44570,
1122 => 44560,
1123 => 44550,
1124 => 44540,
1125 => 44530,
1126 => 44520,
1127 => 44509,
1128 => 44499,
1129 => 44488,
1130 => 44478,
1131 => 44467,
1132 => 44456,
1133 => 44445,
1134 => 44434,
1135 => 44423,
1136 => 44412,
1137 => 44401,
1138 => 44389,
1139 => 44378,
1140 => 44366,
1141 => 44354,
1142 => 44343,
1143 => 44331,
1144 => 44319,
1145 => 44306,
1146 => 44294,
1147 => 44282,
1148 => 44269,
1149 => 44257,
1150 => 44244,
1151 => 44232,
1152 => 44219,
1153 => 44206,
1154 => 44193,
1155 => 44180,
1156 => 44167,
1157 => 44153,
1158 => 44140,
1159 => 44126,
1160 => 44113,
1161 => 44099,
1162 => 44085,
1163 => 44071,
1164 => 44057,
1165 => 44043,
1166 => 44029,
1167 => 44015,
1168 => 44000,
1169 => 43986,
1170 => 43971,
1171 => 43956,
1172 => 43942,
1173 => 43927,
1174 => 43912,
1175 => 43897,
1176 => 43881,
1177 => 43866,
1178 => 43851,
1179 => 43835,
1180 => 43820,
1181 => 43804,
1182 => 43788,
1183 => 43772,
1184 => 43756,
1185 => 43740,
1186 => 43724,
1187 => 43708,
1188 => 43692,
1189 => 43675,
1190 => 43658,
1191 => 43642,
1192 => 43625,
1193 => 43608,
1194 => 43591,
1195 => 43574,
1196 => 43557,
1197 => 43540,
1198 => 43522,
1199 => 43505,
1200 => 43487,
1201 => 43470,
1202 => 43452,
1203 => 43434,
1204 => 43416,
1205 => 43398,
1206 => 43380,
1207 => 43362,
1208 => 43344,
1209 => 43325,
1210 => 43307,
1211 => 43288,
1212 => 43269,
1213 => 43251,
1214 => 43232,
1215 => 43213,
1216 => 43194,
1217 => 43174,
1218 => 43155,
1219 => 43136,
1220 => 43116,
1221 => 43097,
1222 => 43077,
1223 => 43057,
1224 => 43037,
1225 => 43017,
1226 => 42997,
1227 => 42977,
1228 => 42957,
1229 => 42936,
1230 => 42916,
1231 => 42895,
1232 => 42875,
1233 => 42854,
1234 => 42833,
1235 => 42812,
1236 => 42791,
1237 => 42770,
1238 => 42749,
1239 => 42728,
1240 => 42706,
1241 => 42685,
1242 => 42663,
1243 => 42641,
1244 => 42620,
1245 => 42598,
1246 => 42576,
1247 => 42554,
1248 => 42532,
1249 => 42509,
1250 => 42487,
1251 => 42464,
1252 => 42442,
1253 => 42419,
1254 => 42397,
1255 => 42374,
1256 => 42351,
1257 => 42328,
1258 => 42305,
1259 => 42281,
1260 => 42258,
1261 => 42235,
1262 => 42211,
1263 => 42188,
1264 => 42164,
1265 => 42140,
1266 => 42116,
1267 => 42092,
1268 => 42068,
1269 => 42044,
1270 => 42020,
1271 => 41995,
1272 => 41971,
1273 => 41946,
1274 => 41922,
1275 => 41897,
1276 => 41872,
1277 => 41847,
1278 => 41822,
1279 => 41797,
1280 => 41772,
1281 => 41747,
1282 => 41721,
1283 => 41696,
1284 => 41670,
1285 => 41645,
1286 => 41619,
1287 => 41593,
1288 => 41567,
1289 => 41541,
1290 => 41515,
1291 => 41489,
1292 => 41462,
1293 => 41436,
1294 => 41410,
1295 => 41383,
1296 => 41356,
1297 => 41329,
1298 => 41303,
1299 => 41276,
1300 => 41249,
1301 => 41221,
1302 => 41194,
1303 => 41167,
1304 => 41139,
1305 => 41112,
1306 => 41084,
1307 => 41057,
1308 => 41029,
1309 => 41001,
1310 => 40973,
1311 => 40945,
1312 => 40917,
1313 => 40889,
1314 => 40860,
1315 => 40832,
1316 => 40803,
1317 => 40775,
1318 => 40746,
1319 => 40717,
1320 => 40688,
1321 => 40659,
1322 => 40630,
1323 => 40601,
1324 => 40572,
1325 => 40542,
1326 => 40513,
1327 => 40484,
1328 => 40454,
1329 => 40424,
1330 => 40394,
1331 => 40365,
1332 => 40335,
1333 => 40305,
1334 => 40274,
1335 => 40244,
1336 => 40214,
1337 => 40183,
1338 => 40153,
1339 => 40122,
1340 => 40092,
1341 => 40061,
1342 => 40030,
1343 => 39999,
1344 => 39968,
1345 => 39937,
1346 => 39906,
1347 => 39874,
1348 => 39843,
1349 => 39811,
1350 => 39780,
1351 => 39748,
1352 => 39716,
1353 => 39684,
1354 => 39653,
1355 => 39621,
1356 => 39588,
1357 => 39556,
1358 => 39524,
1359 => 39492,
1360 => 39459,
1361 => 39427,
1362 => 39394,
1363 => 39361,
1364 => 39328,
1365 => 39295,
1366 => 39262,
1367 => 39229,
1368 => 39196,
1369 => 39163,
1370 => 39130,
1371 => 39096,
1372 => 39063,
1373 => 39029,
1374 => 38995,
1375 => 38962,
1376 => 38928,
1377 => 38894,
1378 => 38860,
1379 => 38826,
1380 => 38791,
1381 => 38757,
1382 => 38723,
1383 => 38688,
1384 => 38654,
1385 => 38619,
1386 => 38584,
1387 => 38549,
1388 => 38515,
1389 => 38480,
1390 => 38444,
1391 => 38409,
1392 => 38374,
1393 => 38339,
1394 => 38303,
1395 => 38268,
1396 => 38232,
1397 => 38197,
1398 => 38161,
1399 => 38125,
1400 => 38089,
1401 => 38053,
1402 => 38017,
1403 => 37981,
1404 => 37945,
1405 => 37908,
1406 => 37872,
1407 => 37835,
1408 => 37799,
1409 => 37762,
1410 => 37725,
1411 => 37688,
1412 => 37651,
1413 => 37614,
1414 => 37577,
1415 => 37540,
1416 => 37503,
1417 => 37465,
1418 => 37428,
1419 => 37390,
1420 => 37353,
1421 => 37315,
1422 => 37277,
1423 => 37240,
1424 => 37202,
1425 => 37164,
1426 => 37125,
1427 => 37087,
1428 => 37049,
1429 => 37011,
1430 => 36972,
1431 => 36934,
1432 => 36895,
1433 => 36856,
1434 => 36818,
1435 => 36779,
1436 => 36740,
1437 => 36701,
1438 => 36662,
1439 => 36623,
1440 => 36583,
1441 => 36544,
1442 => 36505,
1443 => 36465,
1444 => 36426,
1445 => 36386,
1446 => 36346,
1447 => 36306,
1448 => 36266,
1449 => 36227,
1450 => 36186,
1451 => 36146,
1452 => 36106,
1453 => 36066,
1454 => 36025,
1455 => 35985,
1456 => 35944,
1457 => 35904,
1458 => 35863,
1459 => 35822,
1460 => 35781,
1461 => 35741,
1462 => 35700,
1463 => 35658,
1464 => 35617,
1465 => 35576,
1466 => 35535,
1467 => 35493,
1468 => 35452,
1469 => 35410,
1470 => 35369,
1471 => 35327,
1472 => 35285,
1473 => 35243,
1474 => 35201,
1475 => 35159,
1476 => 35117,
1477 => 35075,
1478 => 35033,
1479 => 34990,
1480 => 34948,
1481 => 34905,
1482 => 34863,
1483 => 34820,
1484 => 34777,
1485 => 34734,
1486 => 34692,
1487 => 34649,
1488 => 34606,
1489 => 34562,
1490 => 34519,
1491 => 34476,
1492 => 34433,
1493 => 34389,
1494 => 34346,
1495 => 34302,
1496 => 34258,
1497 => 34215,
1498 => 34171,
1499 => 34127,
1500 => 34083,
1501 => 34039,
1502 => 33995,
1503 => 33951,
1504 => 33907,
1505 => 33862,
1506 => 33818,
1507 => 33773,
1508 => 33729,
1509 => 33684,
1510 => 33639,
1511 => 33595,
1512 => 33550,
1513 => 33505,
1514 => 33460,
1515 => 33415,
1516 => 33370,
1517 => 33324,
1518 => 33279,
1519 => 33234,
1520 => 33188,
1521 => 33143,
1522 => 33097,
1523 => 33052,
1524 => 33006,
1525 => 32960,
1526 => 32914,
1527 => 32868,
1528 => 32822,
1529 => 32776,
1530 => 32730,
1531 => 32684,
1532 => 32637,
1533 => 32591,
1534 => 32544,
1535 => 32498,
1536 => 32451,
1537 => 32405,
1538 => 32358,
1539 => 32311,
1540 => 32264,
1541 => 32217,
1542 => 32170,
1543 => 32123,
1544 => 32076,
1545 => 32029,
1546 => 31981,
1547 => 31934,
1548 => 31887,
1549 => 31839,
1550 => 31791,
1551 => 31744,
1552 => 31696,
1553 => 31648,
1554 => 31600,
1555 => 31552,
1556 => 31504,
1557 => 31456,
1558 => 31408,
1559 => 31360,
1560 => 31312,
1561 => 31263,
1562 => 31215,
1563 => 31166,
1564 => 31118,
1565 => 31069,
1566 => 31020,
1567 => 30972,
1568 => 30923,
1569 => 30874,
1570 => 30825,
1571 => 30776,
1572 => 30727,
1573 => 30678,
1574 => 30628,
1575 => 30579,
1576 => 30530,
1577 => 30480,
1578 => 30431,
1579 => 30381,
1580 => 30332,
1581 => 30282,
1582 => 30232,
1583 => 30182,
1584 => 30132,
1585 => 30082,
1586 => 30032,
1587 => 29982,
1588 => 29932,
1589 => 29882,
1590 => 29831,
1591 => 29781,
1592 => 29731,
1593 => 29680,
1594 => 29630,
1595 => 29579,
1596 => 29528,
1597 => 29477,
1598 => 29427,
1599 => 29376,
1600 => 29325,
1601 => 29274,
1602 => 29223,
1603 => 29172,
1604 => 29120,
1605 => 29069,
1606 => 29018,
1607 => 28966,
1608 => 28915,
1609 => 28863,
1610 => 28812,
1611 => 28760,
1612 => 28708,
1613 => 28657,
1614 => 28605,
1615 => 28553,
1616 => 28501,
1617 => 28449,
1618 => 28397,
1619 => 28345,
1620 => 28292,
1621 => 28240,
1622 => 28188,
1623 => 28135,
1624 => 28083,
1625 => 28030,
1626 => 27978,
1627 => 27925,
1628 => 27873,
1629 => 27820,
1630 => 27767,
1631 => 27714,
1632 => 27661,
1633 => 27608,
1634 => 27555,
1635 => 27502,
1636 => 27449,
1637 => 27395,
1638 => 27342,
1639 => 27289,
1640 => 27235,
1641 => 27182,
1642 => 27128,
1643 => 27075,
1644 => 27021,
1645 => 26967,
1646 => 26914,
1647 => 26860,
1648 => 26806,
1649 => 26752,
1650 => 26698,
1651 => 26644,
1652 => 26590,
1653 => 26535,
1654 => 26481,
1655 => 26427,
1656 => 26373,
1657 => 26318,
1658 => 26264,
1659 => 26209,
1660 => 26155,
1661 => 26100,
1662 => 26045,
1663 => 25990,
1664 => 25936,
1665 => 25881,
1666 => 25826,
1667 => 25771,
1668 => 25716,
1669 => 25661,
1670 => 25606,
1671 => 25550,
1672 => 25495,
1673 => 25440,
1674 => 25384,
1675 => 25329,
1676 => 25274,
1677 => 25218,
1678 => 25162,
1679 => 25107,
1680 => 25051,
1681 => 24995,
1682 => 24940,
1683 => 24884,
1684 => 24828,
1685 => 24772,
1686 => 24716,
1687 => 24660,
1688 => 24604,
1689 => 24547,
1690 => 24491,
1691 => 24435,
1692 => 24379,
1693 => 24322,
1694 => 24266,
1695 => 24209,
1696 => 24153,
1697 => 24096,
1698 => 24039,
1699 => 23983,
1700 => 23926,
1701 => 23869,
1702 => 23812,
1703 => 23755,
1704 => 23698,
1705 => 23641,
1706 => 23584,
1707 => 23527,
1708 => 23470,
1709 => 23413,
1710 => 23356,
1711 => 23298,
1712 => 23241,
1713 => 23183,
1714 => 23126,
1715 => 23069,
1716 => 23011,
1717 => 22953,
1718 => 22896,
1719 => 22838,
1720 => 22780,
1721 => 22722,
1722 => 22665,
1723 => 22607,
1724 => 22549,
1725 => 22491,
1726 => 22433,
1727 => 22375,
1728 => 22316,
1729 => 22258,
1730 => 22200,
1731 => 22142,
1732 => 22083,
1733 => 22025,
1734 => 21967,
1735 => 21908,
1736 => 21850,
1737 => 21791,
1738 => 21732,
1739 => 21674,
1740 => 21615,
1741 => 21556,
1742 => 21497,
1743 => 21439,
1744 => 21380,
1745 => 21321,
1746 => 21262,
1747 => 21203,
1748 => 21144,
1749 => 21085,
1750 => 21025,
1751 => 20966,
1752 => 20907,
1753 => 20848,
1754 => 20788,
1755 => 20729,
1756 => 20669,
1757 => 20610,
1758 => 20550,
1759 => 20491,
1760 => 20431,
1761 => 20372,
1762 => 20312,
1763 => 20252,
1764 => 20192,
1765 => 20133,
1766 => 20073,
1767 => 20013,
1768 => 19953,
1769 => 19893,
1770 => 19833,
1771 => 19773,
1772 => 19713,
1773 => 19653,
1774 => 19592,
1775 => 19532,
1776 => 19472,
1777 => 19412,
1778 => 19351,
1779 => 19291,
1780 => 19230,
1781 => 19170,
1782 => 19109,
1783 => 19049,
1784 => 18988,
1785 => 18928,
1786 => 18867,
1787 => 18806,
1788 => 18745,
1789 => 18685,
1790 => 18624,
1791 => 18563,
1792 => 18502,
1793 => 18441,
1794 => 18380,
1795 => 18319,
1796 => 18258,
1797 => 18197,
1798 => 18136,
1799 => 18074,
1800 => 18013,
1801 => 17952,
1802 => 17891,
1803 => 17829,
1804 => 17768,
1805 => 17707,
1806 => 17645,
1807 => 17584,
1808 => 17522,
1809 => 17461,
1810 => 17399,
1811 => 17337,
1812 => 17276,
1813 => 17214,
1814 => 17152,
1815 => 17090,
1816 => 17029,
1817 => 16967,
1818 => 16905,
1819 => 16843,
1820 => 16781,
1821 => 16719,
1822 => 16657,
1823 => 16595,
1824 => 16533,
1825 => 16471,
1826 => 16409,
1827 => 16346,
1828 => 16284,
1829 => 16222,
1830 => 16160,
1831 => 16097,
1832 => 16035,
1833 => 15973,
1834 => 15910,
1835 => 15848,
1836 => 15785,
1837 => 15723,
1838 => 15660,
1839 => 15598,
1840 => 15535,
1841 => 15472,
1842 => 15410,
1843 => 15347,
1844 => 15284,
1845 => 15221,
1846 => 15159,
1847 => 15096,
1848 => 15033,
1849 => 14970,
1850 => 14907,
1851 => 14844,
1852 => 14781,
1853 => 14718,
1854 => 14655,
1855 => 14592,
1856 => 14529,
1857 => 14466,
1858 => 14403,
1859 => 14340,
1860 => 14276,
1861 => 14213,
1862 => 14150,
1863 => 14086,
1864 => 14023,
1865 => 13960,
1866 => 13896,
1867 => 13833,
1868 => 13770,
1869 => 13706,
1870 => 13643,
1871 => 13579,
1872 => 13515,
1873 => 13452,
1874 => 13388,
1875 => 13325,
1876 => 13261,
1877 => 13197,
1878 => 13134,
1879 => 13070,
1880 => 13006,
1881 => 12942,
1882 => 12878,
1883 => 12815,
1884 => 12751,
1885 => 12687,
1886 => 12623,
1887 => 12559,
1888 => 12495,
1889 => 12431,
1890 => 12367,
1891 => 12303,
1892 => 12239,
1893 => 12175,
1894 => 12111,
1895 => 12047,
1896 => 11982,
1897 => 11918,
1898 => 11854,
1899 => 11790,
1900 => 11726,
1901 => 11661,
1902 => 11597,
1903 => 11533,
1904 => 11468,
1905 => 11404,
1906 => 11340,
1907 => 11275,
1908 => 11211,
1909 => 11146,
1910 => 11082,
1911 => 11017,
1912 => 10953,
1913 => 10888,
1914 => 10824,
1915 => 10759,
1916 => 10694,
1917 => 10630,
1918 => 10565,
1919 => 10501,
1920 => 10436,
1921 => 10371,
1922 => 10306,
1923 => 10242,
1924 => 10177,
1925 => 10112,
1926 => 10047,
1927 => 9983,
1928 => 9918,
1929 => 9853,
1930 => 9788,
1931 => 9723,
1932 => 9658,
1933 => 9593,
1934 => 9528,
1935 => 9463,
1936 => 9398,
1937 => 9333,
1938 => 9268,
1939 => 9203,
1940 => 9138,
1941 => 9073,
1942 => 9008,
1943 => 8943,
1944 => 8878,
1945 => 8813,
1946 => 8748,
1947 => 8683,
1948 => 8617,
1949 => 8552,
1950 => 8487,
1951 => 8422,
1952 => 8357,
1953 => 8291,
1954 => 8226,
1955 => 8161,
1956 => 8095,
1957 => 8030,
1958 => 7965,
1959 => 7899,
1960 => 7834,
1961 => 7769,
1962 => 7703,
1963 => 7638,
1964 => 7573,
1965 => 7507,
1966 => 7442,
1967 => 7376,
1968 => 7311,
1969 => 7245,
1970 => 7180,
1971 => 7114,
1972 => 7049,
1973 => 6983,
1974 => 6918,
1975 => 6852,
1976 => 6787,
1977 => 6721,
1978 => 6656,
1979 => 6590,
1980 => 6524,
1981 => 6459,
1982 => 6393,
1983 => 6328,
1984 => 6262,
1985 => 6196,
1986 => 6131,
1987 => 6065,
1988 => 5999,
1989 => 5934,
1990 => 5868,
1991 => 5802,
1992 => 5737,
1993 => 5671,
1994 => 5605,
1995 => 5539,
1996 => 5474,
1997 => 5408,
1998 => 5342,
1999 => 5276,
2000 => 5211,
2001 => 5145,
2002 => 5079,
2003 => 5013,
2004 => 4947,
2005 => 4882,
2006 => 4816,
2007 => 4750,
2008 => 4684,
2009 => 4618,
2010 => 4552,
2011 => 4487,
2012 => 4421,
2013 => 4355,
2014 => 4289,
2015 => 4223,
2016 => 4157,
2017 => 4091,
2018 => 4026,
2019 => 3960,
2020 => 3894,
2021 => 3828,
2022 => 3762,
2023 => 3696,
2024 => 3630,
2025 => 3564,
2026 => 3498,
2027 => 3432,
2028 => 3366,
2029 => 3301,
2030 => 3235,
2031 => 3169,
2032 => 3103,
2033 => 3037,
2034 => 2971,
2035 => 2905,
2036 => 2839,
2037 => 2773,
2038 => 2707,
2039 => 2641,
2040 => 2575,
2041 => 2509,
2042 => 2443,
2043 => 2377,
2044 => 2311,
2045 => 2245,
2046 => 2179,
2047 => 2113,
2048 => 2048,
2049 => 1982,
2050 => 1916,
2051 => 1850,
2052 => 1784,
2053 => 1718,
2054 => 1652,
2055 => 1586,
2056 => 1520,
2057 => 1454,
2058 => 1388,
2059 => 1322,
2060 => 1256,
2061 => 1190,
2062 => 1124,
2063 => 1058,
2064 => 992,
2065 => 926,
2066 => 860,
2067 => 794,
2068 => 729,
2069 => 663,
2070 => 597,
2071 => 531,
2072 => 465,
2073 => 399,
2074 => 333,
2075 => 267,
2076 => 201,
2077 => 135,
2078 => 69,
2079 => 4,
2080 => -62,
2081 => -128,
2082 => -194,
2083 => -260,
2084 => -326,
2085 => -392,
2086 => -457,
2087 => -523,
2088 => -589,
2089 => -655,
2090 => -721,
2091 => -787,
2092 => -852,
2093 => -918,
2094 => -984,
2095 => -1050,
2096 => -1116,
2097 => -1181,
2098 => -1247,
2099 => -1313,
2100 => -1379,
2101 => -1444,
2102 => -1510,
2103 => -1576,
2104 => -1642,
2105 => -1707,
2106 => -1773,
2107 => -1839,
2108 => -1904,
2109 => -1970,
2110 => -2036,
2111 => -2101,
2112 => -2167,
2113 => -2233,
2114 => -2298,
2115 => -2364,
2116 => -2429,
2117 => -2495,
2118 => -2561,
2119 => -2626,
2120 => -2692,
2121 => -2757,
2122 => -2823,
2123 => -2888,
2124 => -2954,
2125 => -3019,
2126 => -3085,
2127 => -3150,
2128 => -3216,
2129 => -3281,
2130 => -3347,
2131 => -3412,
2132 => -3478,
2133 => -3543,
2134 => -3608,
2135 => -3674,
2136 => -3739,
2137 => -3804,
2138 => -3870,
2139 => -3935,
2140 => -4000,
2141 => -4066,
2142 => -4131,
2143 => -4196,
2144 => -4262,
2145 => -4327,
2146 => -4392,
2147 => -4457,
2148 => -4522,
2149 => -4588,
2150 => -4653,
2151 => -4718,
2152 => -4783,
2153 => -4848,
2154 => -4913,
2155 => -4978,
2156 => -5043,
2157 => -5108,
2158 => -5173,
2159 => -5238,
2160 => -5303,
2161 => -5368,
2162 => -5433,
2163 => -5498,
2164 => -5563,
2165 => -5628,
2166 => -5693,
2167 => -5758,
2168 => -5823,
2169 => -5888,
2170 => -5952,
2171 => -6017,
2172 => -6082,
2173 => -6147,
2174 => -6211,
2175 => -6276,
2176 => -6341,
2177 => -6406,
2178 => -6470,
2179 => -6535,
2180 => -6599,
2181 => -6664,
2182 => -6729,
2183 => -6793,
2184 => -6858,
2185 => -6922,
2186 => -6987,
2187 => -7051,
2188 => -7116,
2189 => -7180,
2190 => -7245,
2191 => -7309,
2192 => -7373,
2193 => -7438,
2194 => -7502,
2195 => -7566,
2196 => -7631,
2197 => -7695,
2198 => -7759,
2199 => -7823,
2200 => -7887,
2201 => -7952,
2202 => -8016,
2203 => -8080,
2204 => -8144,
2205 => -8208,
2206 => -8272,
2207 => -8336,
2208 => -8400,
2209 => -8464,
2210 => -8528,
2211 => -8592,
2212 => -8656,
2213 => -8720,
2214 => -8783,
2215 => -8847,
2216 => -8911,
2217 => -8975,
2218 => -9039,
2219 => -9102,
2220 => -9166,
2221 => -9230,
2222 => -9293,
2223 => -9357,
2224 => -9420,
2225 => -9484,
2226 => -9548,
2227 => -9611,
2228 => -9675,
2229 => -9738,
2230 => -9801,
2231 => -9865,
2232 => -9928,
2233 => -9991,
2234 => -10055,
2235 => -10118,
2236 => -10181,
2237 => -10245,
2238 => -10308,
2239 => -10371,
2240 => -10434,
2241 => -10497,
2242 => -10560,
2243 => -10623,
2244 => -10686,
2245 => -10749,
2246 => -10812,
2247 => -10875,
2248 => -10938,
2249 => -11001,
2250 => -11064,
2251 => -11126,
2252 => -11189,
2253 => -11252,
2254 => -11315,
2255 => -11377,
2256 => -11440,
2257 => -11503,
2258 => -11565,
2259 => -11628,
2260 => -11690,
2261 => -11753,
2262 => -11815,
2263 => -11878,
2264 => -11940,
2265 => -12002,
2266 => -12065,
2267 => -12127,
2268 => -12189,
2269 => -12251,
2270 => -12314,
2271 => -12376,
2272 => -12438,
2273 => -12500,
2274 => -12562,
2275 => -12624,
2276 => -12686,
2277 => -12748,
2278 => -12810,
2279 => -12872,
2280 => -12934,
2281 => -12995,
2282 => -13057,
2283 => -13119,
2284 => -13181,
2285 => -13242,
2286 => -13304,
2287 => -13366,
2288 => -13427,
2289 => -13489,
2290 => -13550,
2291 => -13612,
2292 => -13673,
2293 => -13734,
2294 => -13796,
2295 => -13857,
2296 => -13918,
2297 => -13979,
2298 => -14041,
2299 => -14102,
2300 => -14163,
2301 => -14224,
2302 => -14285,
2303 => -14346,
2304 => -14407,
2305 => -14468,
2306 => -14529,
2307 => -14590,
2308 => -14650,
2309 => -14711,
2310 => -14772,
2311 => -14833,
2312 => -14893,
2313 => -14954,
2314 => -15014,
2315 => -15075,
2316 => -15135,
2317 => -15196,
2318 => -15256,
2319 => -15317,
2320 => -15377,
2321 => -15437,
2322 => -15497,
2323 => -15558,
2324 => -15618,
2325 => -15678,
2326 => -15738,
2327 => -15798,
2328 => -15858,
2329 => -15918,
2330 => -15978,
2331 => -16038,
2332 => -16097,
2333 => -16157,
2334 => -16217,
2335 => -16277,
2336 => -16336,
2337 => -16396,
2338 => -16455,
2339 => -16515,
2340 => -16574,
2341 => -16634,
2342 => -16693,
2343 => -16753,
2344 => -16812,
2345 => -16871,
2346 => -16930,
2347 => -16990,
2348 => -17049,
2349 => -17108,
2350 => -17167,
2351 => -17226,
2352 => -17285,
2353 => -17344,
2354 => -17402,
2355 => -17461,
2356 => -17520,
2357 => -17579,
2358 => -17637,
2359 => -17696,
2360 => -17755,
2361 => -17813,
2362 => -17872,
2363 => -17930,
2364 => -17988,
2365 => -18047,
2366 => -18105,
2367 => -18163,
2368 => -18221,
2369 => -18280,
2370 => -18338,
2371 => -18396,
2372 => -18454,
2373 => -18512,
2374 => -18570,
2375 => -18627,
2376 => -18685,
2377 => -18743,
2378 => -18801,
2379 => -18858,
2380 => -18916,
2381 => -18974,
2382 => -19031,
2383 => -19088,
2384 => -19146,
2385 => -19203,
2386 => -19261,
2387 => -19318,
2388 => -19375,
2389 => -19432,
2390 => -19489,
2391 => -19546,
2392 => -19603,
2393 => -19660,
2394 => -19717,
2395 => -19774,
2396 => -19831,
2397 => -19888,
2398 => -19944,
2399 => -20001,
2400 => -20058,
2401 => -20114,
2402 => -20171,
2403 => -20227,
2404 => -20284,
2405 => -20340,
2406 => -20396,
2407 => -20452,
2408 => -20509,
2409 => -20565,
2410 => -20621,
2411 => -20677,
2412 => -20733,
2413 => -20789,
2414 => -20845,
2415 => -20900,
2416 => -20956,
2417 => -21012,
2418 => -21067,
2419 => -21123,
2420 => -21179,
2421 => -21234,
2422 => -21289,
2423 => -21345,
2424 => -21400,
2425 => -21455,
2426 => -21511,
2427 => -21566,
2428 => -21621,
2429 => -21676,
2430 => -21731,
2431 => -21786,
2432 => -21841,
2433 => -21895,
2434 => -21950,
2435 => -22005,
2436 => -22060,
2437 => -22114,
2438 => -22169,
2439 => -22223,
2440 => -22278,
2441 => -22332,
2442 => -22386,
2443 => -22440,
2444 => -22495,
2445 => -22549,
2446 => -22603,
2447 => -22657,
2448 => -22711,
2449 => -22765,
2450 => -22819,
2451 => -22872,
2452 => -22926,
2453 => -22980,
2454 => -23033,
2455 => -23087,
2456 => -23140,
2457 => -23194,
2458 => -23247,
2459 => -23300,
2460 => -23354,
2461 => -23407,
2462 => -23460,
2463 => -23513,
2464 => -23566,
2465 => -23619,
2466 => -23672,
2467 => -23725,
2468 => -23778,
2469 => -23830,
2470 => -23883,
2471 => -23935,
2472 => -23988,
2473 => -24040,
2474 => -24093,
2475 => -24145,
2476 => -24197,
2477 => -24250,
2478 => -24302,
2479 => -24354,
2480 => -24406,
2481 => -24458,
2482 => -24510,
2483 => -24562,
2484 => -24613,
2485 => -24665,
2486 => -24717,
2487 => -24768,
2488 => -24820,
2489 => -24871,
2490 => -24923,
2491 => -24974,
2492 => -25025,
2493 => -25077,
2494 => -25128,
2495 => -25179,
2496 => -25230,
2497 => -25281,
2498 => -25332,
2499 => -25382,
2500 => -25433,
2501 => -25484,
2502 => -25535,
2503 => -25585,
2504 => -25636,
2505 => -25686,
2506 => -25736,
2507 => -25787,
2508 => -25837,
2509 => -25887,
2510 => -25937,
2511 => -25987,
2512 => -26037,
2513 => -26087,
2514 => -26137,
2515 => -26187,
2516 => -26237,
2517 => -26286,
2518 => -26336,
2519 => -26385,
2520 => -26435,
2521 => -26484,
2522 => -26533,
2523 => -26583,
2524 => -26632,
2525 => -26681,
2526 => -26730,
2527 => -26779,
2528 => -26828,
2529 => -26877,
2530 => -26925,
2531 => -26974,
2532 => -27023,
2533 => -27071,
2534 => -27120,
2535 => -27168,
2536 => -27217,
2537 => -27265,
2538 => -27313,
2539 => -27361,
2540 => -27409,
2541 => -27457,
2542 => -27505,
2543 => -27553,
2544 => -27601,
2545 => -27649,
2546 => -27696,
2547 => -27744,
2548 => -27792,
2549 => -27839,
2550 => -27886,
2551 => -27934,
2552 => -27981,
2553 => -28028,
2554 => -28075,
2555 => -28122,
2556 => -28169,
2557 => -28216,
2558 => -28263,
2559 => -28310,
2560 => -28356,
2561 => -28403,
2562 => -28449,
2563 => -28496,
2564 => -28542,
2565 => -28589,
2566 => -28635,
2567 => -28681,
2568 => -28727,
2569 => -28773,
2570 => -28819,
2571 => -28865,
2572 => -28911,
2573 => -28957,
2574 => -29002,
2575 => -29048,
2576 => -29093,
2577 => -29139,
2578 => -29184,
2579 => -29229,
2580 => -29275,
2581 => -29320,
2582 => -29365,
2583 => -29410,
2584 => -29455,
2585 => -29500,
2586 => -29544,
2587 => -29589,
2588 => -29634,
2589 => -29678,
2590 => -29723,
2591 => -29767,
2592 => -29812,
2593 => -29856,
2594 => -29900,
2595 => -29944,
2596 => -29988,
2597 => -30032,
2598 => -30076,
2599 => -30120,
2600 => -30163,
2601 => -30207,
2602 => -30251,
2603 => -30294,
2604 => -30338,
2605 => -30381,
2606 => -30424,
2607 => -30467,
2608 => -30511,
2609 => -30554,
2610 => -30597,
2611 => -30639,
2612 => -30682,
2613 => -30725,
2614 => -30768,
2615 => -30810,
2616 => -30853,
2617 => -30895,
2618 => -30938,
2619 => -30980,
2620 => -31022,
2621 => -31064,
2622 => -31106,
2623 => -31148,
2624 => -31190,
2625 => -31232,
2626 => -31274,
2627 => -31315,
2628 => -31357,
2629 => -31398,
2630 => -31440,
2631 => -31481,
2632 => -31522,
2633 => -31563,
2634 => -31605,
2635 => -31646,
2636 => -31686,
2637 => -31727,
2638 => -31768,
2639 => -31809,
2640 => -31849,
2641 => -31890,
2642 => -31930,
2643 => -31971,
2644 => -32011,
2645 => -32051,
2646 => -32091,
2647 => -32132,
2648 => -32171,
2649 => -32211,
2650 => -32251,
2651 => -32291,
2652 => -32331,
2653 => -32370,
2654 => -32410,
2655 => -32449,
2656 => -32488,
2657 => -32528,
2658 => -32567,
2659 => -32606,
2660 => -32645,
2661 => -32684,
2662 => -32723,
2663 => -32761,
2664 => -32800,
2665 => -32839,
2666 => -32877,
2667 => -32916,
2668 => -32954,
2669 => -32992,
2670 => -33030,
2671 => -33069,
2672 => -33107,
2673 => -33145,
2674 => -33182,
2675 => -33220,
2676 => -33258,
2677 => -33295,
2678 => -33333,
2679 => -33370,
2680 => -33408,
2681 => -33445,
2682 => -33482,
2683 => -33519,
2684 => -33556,
2685 => -33593,
2686 => -33630,
2687 => -33667,
2688 => -33704,
2689 => -33740,
2690 => -33777,
2691 => -33813,
2692 => -33850,
2693 => -33886,
2694 => -33922,
2695 => -33958,
2696 => -33994,
2697 => -34030,
2698 => -34066,
2699 => -34102,
2700 => -34137,
2701 => -34173,
2702 => -34208,
2703 => -34244,
2704 => -34279,
2705 => -34314,
2706 => -34349,
2707 => -34385,
2708 => -34420,
2709 => -34454,
2710 => -34489,
2711 => -34524,
2712 => -34559,
2713 => -34593,
2714 => -34628,
2715 => -34662,
2716 => -34696,
2717 => -34731,
2718 => -34765,
2719 => -34799,
2720 => -34833,
2721 => -34867,
2722 => -34900,
2723 => -34934,
2724 => -34968,
2725 => -35001,
2726 => -35035,
2727 => -35068,
2728 => -35101,
2729 => -35134,
2730 => -35167,
2731 => -35200,
2732 => -35233,
2733 => -35266,
2734 => -35299,
2735 => -35332,
2736 => -35364,
2737 => -35397,
2738 => -35429,
2739 => -35461,
2740 => -35493,
2741 => -35526,
2742 => -35558,
2743 => -35589,
2744 => -35621,
2745 => -35653,
2746 => -35685,
2747 => -35716,
2748 => -35748,
2749 => -35779,
2750 => -35811,
2751 => -35842,
2752 => -35873,
2753 => -35904,
2754 => -35935,
2755 => -35966,
2756 => -35997,
2757 => -36027,
2758 => -36058,
2759 => -36088,
2760 => -36119,
2761 => -36149,
2762 => -36179,
2763 => -36210,
2764 => -36240,
2765 => -36270,
2766 => -36299,
2767 => -36329,
2768 => -36359,
2769 => -36389,
2770 => -36418,
2771 => -36447,
2772 => -36477,
2773 => -36506,
2774 => -36535,
2775 => -36564,
2776 => -36593,
2777 => -36622,
2778 => -36651,
2779 => -36680,
2780 => -36708,
2781 => -36737,
2782 => -36765,
2783 => -36794,
2784 => -36822,
2785 => -36850,
2786 => -36878,
2787 => -36906,
2788 => -36934,
2789 => -36962,
2790 => -36989,
2791 => -37017,
2792 => -37044,
2793 => -37072,
2794 => -37099,
2795 => -37126,
2796 => -37154,
2797 => -37181,
2798 => -37208,
2799 => -37234,
2800 => -37261,
2801 => -37288,
2802 => -37315,
2803 => -37341,
2804 => -37367,
2805 => -37394,
2806 => -37420,
2807 => -37446,
2808 => -37472,
2809 => -37498,
2810 => -37524,
2811 => -37550,
2812 => -37575,
2813 => -37601,
2814 => -37626,
2815 => -37652,
2816 => -37677,
2817 => -37702,
2818 => -37727,
2819 => -37752,
2820 => -37777,
2821 => -37802,
2822 => -37827,
2823 => -37851,
2824 => -37876,
2825 => -37900,
2826 => -37925,
2827 => -37949,
2828 => -37973,
2829 => -37997,
2830 => -38021,
2831 => -38045,
2832 => -38069,
2833 => -38093,
2834 => -38116,
2835 => -38140,
2836 => -38163,
2837 => -38186,
2838 => -38210,
2839 => -38233,
2840 => -38256,
2841 => -38279,
2842 => -38302,
2843 => -38324,
2844 => -38347,
2845 => -38369,
2846 => -38392,
2847 => -38414,
2848 => -38437,
2849 => -38459,
2850 => -38481,
2851 => -38503,
2852 => -38525,
2853 => -38546,
2854 => -38568,
2855 => -38590,
2856 => -38611,
2857 => -38633,
2858 => -38654,
2859 => -38675,
2860 => -38696,
2861 => -38717,
2862 => -38738,
2863 => -38759,
2864 => -38780,
2865 => -38800,
2866 => -38821,
2867 => -38841,
2868 => -38862,
2869 => -38882,
2870 => -38902,
2871 => -38922,
2872 => -38942,
2873 => -38962,
2874 => -38982,
2875 => -39002,
2876 => -39021,
2877 => -39041,
2878 => -39060,
2879 => -39079,
2880 => -39099,
2881 => -39118,
2882 => -39137,
2883 => -39156,
2884 => -39174,
2885 => -39193,
2886 => -39212,
2887 => -39230,
2888 => -39249,
2889 => -39267,
2890 => -39285,
2891 => -39303,
2892 => -39321,
2893 => -39339,
2894 => -39357,
2895 => -39375,
2896 => -39392,
2897 => -39410,
2898 => -39427,
2899 => -39445,
2900 => -39462,
2901 => -39479,
2902 => -39496,
2903 => -39513,
2904 => -39530,
2905 => -39547,
2906 => -39563,
2907 => -39580,
2908 => -39597,
2909 => -39613,
2910 => -39629,
2911 => -39645,
2912 => -39661,
2913 => -39677,
2914 => -39693,
2915 => -39709,
2916 => -39725,
2917 => -39740,
2918 => -39756,
2919 => -39771,
2920 => -39786,
2921 => -39802,
2922 => -39817,
2923 => -39832,
2924 => -39847,
2925 => -39861,
2926 => -39876,
2927 => -39891,
2928 => -39905,
2929 => -39920,
2930 => -39934,
2931 => -39948,
2932 => -39962,
2933 => -39976,
2934 => -39990,
2935 => -40004,
2936 => -40018,
2937 => -40031,
2938 => -40045,
2939 => -40058,
2940 => -40072,
2941 => -40085,
2942 => -40098,
2943 => -40111,
2944 => -40124,
2945 => -40137,
2946 => -40149,
2947 => -40162,
2948 => -40174,
2949 => -40187,
2950 => -40199,
2951 => -40211,
2952 => -40224,
2953 => -40236,
2954 => -40248,
2955 => -40259,
2956 => -40271,
2957 => -40283,
2958 => -40294,
2959 => -40306,
2960 => -40317,
2961 => -40328,
2962 => -40339,
2963 => -40350,
2964 => -40361,
2965 => -40372,
2966 => -40383,
2967 => -40393,
2968 => -40404,
2969 => -40414,
2970 => -40425,
2971 => -40435,
2972 => -40445,
2973 => -40455,
2974 => -40465,
2975 => -40475,
2976 => -40485,
2977 => -40494,
2978 => -40504,
2979 => -40513,
2980 => -40523,
2981 => -40532,
2982 => -40541,
2983 => -40550,
2984 => -40559,
2985 => -40568,
2986 => -40576,
2987 => -40585,
2988 => -40594,
2989 => -40602,
2990 => -40610,
2991 => -40619,
2992 => -40627,
2993 => -40635,
2994 => -40643,
2995 => -40650,
2996 => -40658,
2997 => -40666,
2998 => -40673,
2999 => -40681,
3000 => -40688,
3001 => -40695,
3002 => -40702,
3003 => -40709,
3004 => -40716,
3005 => -40723,
3006 => -40730,
3007 => -40736,
3008 => -40743,
3009 => -40749,
3010 => -40756,
3011 => -40762,
3012 => -40768,
3013 => -40774,
3014 => -40780,
3015 => -40786,
3016 => -40791,
3017 => -40797,
3018 => -40803,
3019 => -40808,
3020 => -40813,
3021 => -40818,
3022 => -40824,
3023 => -40829,
3024 => -40833,
3025 => -40838,
3026 => -40843,
3027 => -40848,
3028 => -40852,
3029 => -40856,
3030 => -40861,
3031 => -40865,
3032 => -40869,
3033 => -40873,
3034 => -40877,
3035 => -40881,
3036 => -40884,
3037 => -40888,
3038 => -40892,
3039 => -40895,
3040 => -40898,
3041 => -40901,
3042 => -40904,
3043 => -40907,
3044 => -40910,
3045 => -40913,
3046 => -40916,
3047 => -40918,
3048 => -40921,
3049 => -40923,
3050 => -40926,
3051 => -40928,
3052 => -40930,
3053 => -40932,
3054 => -40934,
3055 => -40935,
3056 => -40937,
3057 => -40939,
3058 => -40940,
3059 => -40941,
3060 => -40943,
3061 => -40944,
3062 => -40945,
3063 => -40946,
3064 => -40947,
3065 => -40948,
3066 => -40948,
3067 => -40949,
3068 => -40949,
3069 => -40950,
3070 => -40950,
3071 => -40950,
3072 => -40950,
3073 => -40950,
3074 => -40950,
3075 => -40950,
3076 => -40949,
3077 => -40949,
3078 => -40948,
3079 => -40948,
3080 => -40947,
3081 => -40946,
3082 => -40945,
3083 => -40944,
3084 => -40943,
3085 => -40941,
3086 => -40940,
3087 => -40939,
3088 => -40937,
3089 => -40935,
3090 => -40934,
3091 => -40932,
3092 => -40930,
3093 => -40928,
3094 => -40926,
3095 => -40923,
3096 => -40921,
3097 => -40918,
3098 => -40916,
3099 => -40913,
3100 => -40910,
3101 => -40907,
3102 => -40904,
3103 => -40901,
3104 => -40898,
3105 => -40895,
3106 => -40892,
3107 => -40888,
3108 => -40884,
3109 => -40881,
3110 => -40877,
3111 => -40873,
3112 => -40869,
3113 => -40865,
3114 => -40861,
3115 => -40856,
3116 => -40852,
3117 => -40848,
3118 => -40843,
3119 => -40838,
3120 => -40833,
3121 => -40829,
3122 => -40824,
3123 => -40818,
3124 => -40813,
3125 => -40808,
3126 => -40803,
3127 => -40797,
3128 => -40791,
3129 => -40786,
3130 => -40780,
3131 => -40774,
3132 => -40768,
3133 => -40762,
3134 => -40756,
3135 => -40749,
3136 => -40743,
3137 => -40736,
3138 => -40730,
3139 => -40723,
3140 => -40716,
3141 => -40709,
3142 => -40702,
3143 => -40695,
3144 => -40688,
3145 => -40681,
3146 => -40673,
3147 => -40666,
3148 => -40658,
3149 => -40650,
3150 => -40643,
3151 => -40635,
3152 => -40627,
3153 => -40619,
3154 => -40610,
3155 => -40602,
3156 => -40594,
3157 => -40585,
3158 => -40576,
3159 => -40568,
3160 => -40559,
3161 => -40550,
3162 => -40541,
3163 => -40532,
3164 => -40523,
3165 => -40513,
3166 => -40504,
3167 => -40494,
3168 => -40485,
3169 => -40475,
3170 => -40465,
3171 => -40455,
3172 => -40445,
3173 => -40435,
3174 => -40425,
3175 => -40414,
3176 => -40404,
3177 => -40393,
3178 => -40383,
3179 => -40372,
3180 => -40361,
3181 => -40350,
3182 => -40339,
3183 => -40328,
3184 => -40317,
3185 => -40306,
3186 => -40294,
3187 => -40283,
3188 => -40271,
3189 => -40259,
3190 => -40248,
3191 => -40236,
3192 => -40224,
3193 => -40211,
3194 => -40199,
3195 => -40187,
3196 => -40174,
3197 => -40162,
3198 => -40149,
3199 => -40137,
3200 => -40124,
3201 => -40111,
3202 => -40098,
3203 => -40085,
3204 => -40072,
3205 => -40058,
3206 => -40045,
3207 => -40031,
3208 => -40018,
3209 => -40004,
3210 => -39990,
3211 => -39976,
3212 => -39962,
3213 => -39948,
3214 => -39934,
3215 => -39920,
3216 => -39905,
3217 => -39891,
3218 => -39876,
3219 => -39861,
3220 => -39847,
3221 => -39832,
3222 => -39817,
3223 => -39802,
3224 => -39786,
3225 => -39771,
3226 => -39756,
3227 => -39740,
3228 => -39725,
3229 => -39709,
3230 => -39693,
3231 => -39677,
3232 => -39661,
3233 => -39645,
3234 => -39629,
3235 => -39613,
3236 => -39597,
3237 => -39580,
3238 => -39563,
3239 => -39547,
3240 => -39530,
3241 => -39513,
3242 => -39496,
3243 => -39479,
3244 => -39462,
3245 => -39445,
3246 => -39427,
3247 => -39410,
3248 => -39392,
3249 => -39375,
3250 => -39357,
3251 => -39339,
3252 => -39321,
3253 => -39303,
3254 => -39285,
3255 => -39267,
3256 => -39249,
3257 => -39230,
3258 => -39212,
3259 => -39193,
3260 => -39174,
3261 => -39156,
3262 => -39137,
3263 => -39118,
3264 => -39099,
3265 => -39079,
3266 => -39060,
3267 => -39041,
3268 => -39021,
3269 => -39002,
3270 => -38982,
3271 => -38962,
3272 => -38942,
3273 => -38922,
3274 => -38902,
3275 => -38882,
3276 => -38862,
3277 => -38841,
3278 => -38821,
3279 => -38800,
3280 => -38780,
3281 => -38759,
3282 => -38738,
3283 => -38717,
3284 => -38696,
3285 => -38675,
3286 => -38654,
3287 => -38633,
3288 => -38611,
3289 => -38590,
3290 => -38568,
3291 => -38546,
3292 => -38525,
3293 => -38503,
3294 => -38481,
3295 => -38459,
3296 => -38437,
3297 => -38414,
3298 => -38392,
3299 => -38369,
3300 => -38347,
3301 => -38324,
3302 => -38302,
3303 => -38279,
3304 => -38256,
3305 => -38233,
3306 => -38210,
3307 => -38186,
3308 => -38163,
3309 => -38140,
3310 => -38116,
3311 => -38093,
3312 => -38069,
3313 => -38045,
3314 => -38021,
3315 => -37997,
3316 => -37973,
3317 => -37949,
3318 => -37925,
3319 => -37900,
3320 => -37876,
3321 => -37851,
3322 => -37827,
3323 => -37802,
3324 => -37777,
3325 => -37752,
3326 => -37727,
3327 => -37702,
3328 => -37677,
3329 => -37652,
3330 => -37626,
3331 => -37601,
3332 => -37575,
3333 => -37550,
3334 => -37524,
3335 => -37498,
3336 => -37472,
3337 => -37446,
3338 => -37420,
3339 => -37394,
3340 => -37367,
3341 => -37341,
3342 => -37315,
3343 => -37288,
3344 => -37261,
3345 => -37234,
3346 => -37208,
3347 => -37181,
3348 => -37154,
3349 => -37126,
3350 => -37099,
3351 => -37072,
3352 => -37044,
3353 => -37017,
3354 => -36989,
3355 => -36962,
3356 => -36934,
3357 => -36906,
3358 => -36878,
3359 => -36850,
3360 => -36822,
3361 => -36794,
3362 => -36765,
3363 => -36737,
3364 => -36708,
3365 => -36680,
3366 => -36651,
3367 => -36622,
3368 => -36593,
3369 => -36564,
3370 => -36535,
3371 => -36506,
3372 => -36477,
3373 => -36447,
3374 => -36418,
3375 => -36389,
3376 => -36359,
3377 => -36329,
3378 => -36299,
3379 => -36270,
3380 => -36240,
3381 => -36210,
3382 => -36179,
3383 => -36149,
3384 => -36119,
3385 => -36088,
3386 => -36058,
3387 => -36027,
3388 => -35997,
3389 => -35966,
3390 => -35935,
3391 => -35904,
3392 => -35873,
3393 => -35842,
3394 => -35811,
3395 => -35779,
3396 => -35748,
3397 => -35716,
3398 => -35685,
3399 => -35653,
3400 => -35621,
3401 => -35589,
3402 => -35558,
3403 => -35526,
3404 => -35493,
3405 => -35461,
3406 => -35429,
3407 => -35397,
3408 => -35364,
3409 => -35332,
3410 => -35299,
3411 => -35266,
3412 => -35233,
3413 => -35200,
3414 => -35167,
3415 => -35134,
3416 => -35101,
3417 => -35068,
3418 => -35035,
3419 => -35001,
3420 => -34968,
3421 => -34934,
3422 => -34900,
3423 => -34867,
3424 => -34833,
3425 => -34799,
3426 => -34765,
3427 => -34731,
3428 => -34696,
3429 => -34662,
3430 => -34628,
3431 => -34593,
3432 => -34559,
3433 => -34524,
3434 => -34489,
3435 => -34454,
3436 => -34420,
3437 => -34385,
3438 => -34349,
3439 => -34314,
3440 => -34279,
3441 => -34244,
3442 => -34208,
3443 => -34173,
3444 => -34137,
3445 => -34102,
3446 => -34066,
3447 => -34030,
3448 => -33994,
3449 => -33958,
3450 => -33922,
3451 => -33886,
3452 => -33850,
3453 => -33813,
3454 => -33777,
3455 => -33740,
3456 => -33704,
3457 => -33667,
3458 => -33630,
3459 => -33593,
3460 => -33556,
3461 => -33519,
3462 => -33482,
3463 => -33445,
3464 => -33408,
3465 => -33370,
3466 => -33333,
3467 => -33295,
3468 => -33258,
3469 => -33220,
3470 => -33182,
3471 => -33145,
3472 => -33107,
3473 => -33069,
3474 => -33030,
3475 => -32992,
3476 => -32954,
3477 => -32916,
3478 => -32877,
3479 => -32839,
3480 => -32800,
3481 => -32761,
3482 => -32723,
3483 => -32684,
3484 => -32645,
3485 => -32606,
3486 => -32567,
3487 => -32528,
3488 => -32488,
3489 => -32449,
3490 => -32410,
3491 => -32370,
3492 => -32331,
3493 => -32291,
3494 => -32251,
3495 => -32211,
3496 => -32171,
3497 => -32132,
3498 => -32091,
3499 => -32051,
3500 => -32011,
3501 => -31971,
3502 => -31930,
3503 => -31890,
3504 => -31849,
3505 => -31809,
3506 => -31768,
3507 => -31727,
3508 => -31686,
3509 => -31646,
3510 => -31605,
3511 => -31563,
3512 => -31522,
3513 => -31481,
3514 => -31440,
3515 => -31398,
3516 => -31357,
3517 => -31315,
3518 => -31274,
3519 => -31232,
3520 => -31190,
3521 => -31148,
3522 => -31106,
3523 => -31064,
3524 => -31022,
3525 => -30980,
3526 => -30938,
3527 => -30895,
3528 => -30853,
3529 => -30810,
3530 => -30768,
3531 => -30725,
3532 => -30682,
3533 => -30639,
3534 => -30597,
3535 => -30554,
3536 => -30511,
3537 => -30467,
3538 => -30424,
3539 => -30381,
3540 => -30338,
3541 => -30294,
3542 => -30251,
3543 => -30207,
3544 => -30163,
3545 => -30120,
3546 => -30076,
3547 => -30032,
3548 => -29988,
3549 => -29944,
3550 => -29900,
3551 => -29856,
3552 => -29812,
3553 => -29767,
3554 => -29723,
3555 => -29678,
3556 => -29634,
3557 => -29589,
3558 => -29544,
3559 => -29500,
3560 => -29455,
3561 => -29410,
3562 => -29365,
3563 => -29320,
3564 => -29275,
3565 => -29229,
3566 => -29184,
3567 => -29139,
3568 => -29093,
3569 => -29048,
3570 => -29002,
3571 => -28957,
3572 => -28911,
3573 => -28865,
3574 => -28819,
3575 => -28773,
3576 => -28727,
3577 => -28681,
3578 => -28635,
3579 => -28589,
3580 => -28542,
3581 => -28496,
3582 => -28449,
3583 => -28403,
3584 => -28356,
3585 => -28310,
3586 => -28263,
3587 => -28216,
3588 => -28169,
3589 => -28122,
3590 => -28075,
3591 => -28028,
3592 => -27981,
3593 => -27934,
3594 => -27886,
3595 => -27839,
3596 => -27792,
3597 => -27744,
3598 => -27696,
3599 => -27649,
3600 => -27601,
3601 => -27553,
3602 => -27505,
3603 => -27457,
3604 => -27409,
3605 => -27361,
3606 => -27313,
3607 => -27265,
3608 => -27217,
3609 => -27168,
3610 => -27120,
3611 => -27071,
3612 => -27023,
3613 => -26974,
3614 => -26925,
3615 => -26877,
3616 => -26828,
3617 => -26779,
3618 => -26730,
3619 => -26681,
3620 => -26632,
3621 => -26583,
3622 => -26533,
3623 => -26484,
3624 => -26435,
3625 => -26385,
3626 => -26336,
3627 => -26286,
3628 => -26237,
3629 => -26187,
3630 => -26137,
3631 => -26087,
3632 => -26037,
3633 => -25987,
3634 => -25937,
3635 => -25887,
3636 => -25837,
3637 => -25787,
3638 => -25736,
3639 => -25686,
3640 => -25636,
3641 => -25585,
3642 => -25535,
3643 => -25484,
3644 => -25433,
3645 => -25382,
3646 => -25332,
3647 => -25281,
3648 => -25230,
3649 => -25179,
3650 => -25128,
3651 => -25077,
3652 => -25025,
3653 => -24974,
3654 => -24923,
3655 => -24871,
3656 => -24820,
3657 => -24768,
3658 => -24717,
3659 => -24665,
3660 => -24613,
3661 => -24562,
3662 => -24510,
3663 => -24458,
3664 => -24406,
3665 => -24354,
3666 => -24302,
3667 => -24250,
3668 => -24197,
3669 => -24145,
3670 => -24093,
3671 => -24040,
3672 => -23988,
3673 => -23935,
3674 => -23883,
3675 => -23830,
3676 => -23778,
3677 => -23725,
3678 => -23672,
3679 => -23619,
3680 => -23566,
3681 => -23513,
3682 => -23460,
3683 => -23407,
3684 => -23354,
3685 => -23300,
3686 => -23247,
3687 => -23194,
3688 => -23140,
3689 => -23087,
3690 => -23033,
3691 => -22980,
3692 => -22926,
3693 => -22872,
3694 => -22819,
3695 => -22765,
3696 => -22711,
3697 => -22657,
3698 => -22603,
3699 => -22549,
3700 => -22495,
3701 => -22440,
3702 => -22386,
3703 => -22332,
3704 => -22278,
3705 => -22223,
3706 => -22169,
3707 => -22114,
3708 => -22060,
3709 => -22005,
3710 => -21950,
3711 => -21895,
3712 => -21841,
3713 => -21786,
3714 => -21731,
3715 => -21676,
3716 => -21621,
3717 => -21566,
3718 => -21511,
3719 => -21455,
3720 => -21400,
3721 => -21345,
3722 => -21289,
3723 => -21234,
3724 => -21179,
3725 => -21123,
3726 => -21067,
3727 => -21012,
3728 => -20956,
3729 => -20900,
3730 => -20845,
3731 => -20789,
3732 => -20733,
3733 => -20677,
3734 => -20621,
3735 => -20565,
3736 => -20509,
3737 => -20452,
3738 => -20396,
3739 => -20340,
3740 => -20284,
3741 => -20227,
3742 => -20171,
3743 => -20114,
3744 => -20058,
3745 => -20001,
3746 => -19944,
3747 => -19888,
3748 => -19831,
3749 => -19774,
3750 => -19717,
3751 => -19660,
3752 => -19603,
3753 => -19546,
3754 => -19489,
3755 => -19432,
3756 => -19375,
3757 => -19318,
3758 => -19261,
3759 => -19203,
3760 => -19146,
3761 => -19088,
3762 => -19031,
3763 => -18974,
3764 => -18916,
3765 => -18858,
3766 => -18801,
3767 => -18743,
3768 => -18685,
3769 => -18627,
3770 => -18570,
3771 => -18512,
3772 => -18454,
3773 => -18396,
3774 => -18338,
3775 => -18280,
3776 => -18221,
3777 => -18163,
3778 => -18105,
3779 => -18047,
3780 => -17988,
3781 => -17930,
3782 => -17872,
3783 => -17813,
3784 => -17755,
3785 => -17696,
3786 => -17637,
3787 => -17579,
3788 => -17520,
3789 => -17461,
3790 => -17402,
3791 => -17344,
3792 => -17285,
3793 => -17226,
3794 => -17167,
3795 => -17108,
3796 => -17049,
3797 => -16990,
3798 => -16930,
3799 => -16871,
3800 => -16812,
3801 => -16753,
3802 => -16693,
3803 => -16634,
3804 => -16574,
3805 => -16515,
3806 => -16455,
3807 => -16396,
3808 => -16336,
3809 => -16277,
3810 => -16217,
3811 => -16157,
3812 => -16097,
3813 => -16038,
3814 => -15978,
3815 => -15918,
3816 => -15858,
3817 => -15798,
3818 => -15738,
3819 => -15678,
3820 => -15618,
3821 => -15558,
3822 => -15497,
3823 => -15437,
3824 => -15377,
3825 => -15317,
3826 => -15256,
3827 => -15196,
3828 => -15135,
3829 => -15075,
3830 => -15014,
3831 => -14954,
3832 => -14893,
3833 => -14833,
3834 => -14772,
3835 => -14711,
3836 => -14650,
3837 => -14590,
3838 => -14529,
3839 => -14468,
3840 => -14407,
3841 => -14346,
3842 => -14285,
3843 => -14224,
3844 => -14163,
3845 => -14102,
3846 => -14041,
3847 => -13979,
3848 => -13918,
3849 => -13857,
3850 => -13796,
3851 => -13734,
3852 => -13673,
3853 => -13612,
3854 => -13550,
3855 => -13489,
3856 => -13427,
3857 => -13366,
3858 => -13304,
3859 => -13242,
3860 => -13181,
3861 => -13119,
3862 => -13057,
3863 => -12995,
3864 => -12934,
3865 => -12872,
3866 => -12810,
3867 => -12748,
3868 => -12686,
3869 => -12624,
3870 => -12562,
3871 => -12500,
3872 => -12438,
3873 => -12376,
3874 => -12314,
3875 => -12251,
3876 => -12189,
3877 => -12127,
3878 => -12065,
3879 => -12002,
3880 => -11940,
3881 => -11878,
3882 => -11815,
3883 => -11753,
3884 => -11690,
3885 => -11628,
3886 => -11565,
3887 => -11503,
3888 => -11440,
3889 => -11377,
3890 => -11315,
3891 => -11252,
3892 => -11189,
3893 => -11126,
3894 => -11064,
3895 => -11001,
3896 => -10938,
3897 => -10875,
3898 => -10812,
3899 => -10749,
3900 => -10686,
3901 => -10623,
3902 => -10560,
3903 => -10497,
3904 => -10434,
3905 => -10371,
3906 => -10308,
3907 => -10245,
3908 => -10181,
3909 => -10118,
3910 => -10055,
3911 => -9991,
3912 => -9928,
3913 => -9865,
3914 => -9801,
3915 => -9738,
3916 => -9675,
3917 => -9611,
3918 => -9548,
3919 => -9484,
3920 => -9420,
3921 => -9357,
3922 => -9293,
3923 => -9230,
3924 => -9166,
3925 => -9102,
3926 => -9039,
3927 => -8975,
3928 => -8911,
3929 => -8847,
3930 => -8783,
3931 => -8720,
3932 => -8656,
3933 => -8592,
3934 => -8528,
3935 => -8464,
3936 => -8400,
3937 => -8336,
3938 => -8272,
3939 => -8208,
3940 => -8144,
3941 => -8080,
3942 => -8016,
3943 => -7952,
3944 => -7887,
3945 => -7823,
3946 => -7759,
3947 => -7695,
3948 => -7631,
3949 => -7566,
3950 => -7502,
3951 => -7438,
3952 => -7373,
3953 => -7309,
3954 => -7245,
3955 => -7180,
3956 => -7116,
3957 => -7051,
3958 => -6987,
3959 => -6922,
3960 => -6858,
3961 => -6793,
3962 => -6729,
3963 => -6664,
3964 => -6599,
3965 => -6535,
3966 => -6470,
3967 => -6406,
3968 => -6341,
3969 => -6276,
3970 => -6211,
3971 => -6147,
3972 => -6082,
3973 => -6017,
3974 => -5952,
3975 => -5888,
3976 => -5823,
3977 => -5758,
3978 => -5693,
3979 => -5628,
3980 => -5563,
3981 => -5498,
3982 => -5433,
3983 => -5368,
3984 => -5303,
3985 => -5238,
3986 => -5173,
3987 => -5108,
3988 => -5043,
3989 => -4978,
3990 => -4913,
3991 => -4848,
3992 => -4783,
3993 => -4718,
3994 => -4653,
3995 => -4588,
3996 => -4522,
3997 => -4457,
3998 => -4392,
3999 => -4327,
4000 => -4262,
4001 => -4196,
4002 => -4131,
4003 => -4066,
4004 => -4000,
4005 => -3935,
4006 => -3870,
4007 => -3804,
4008 => -3739,
4009 => -3674,
4010 => -3608,
4011 => -3543,
4012 => -3478,
4013 => -3412,
4014 => -3347,
4015 => -3281,
4016 => -3216,
4017 => -3150,
4018 => -3085,
4019 => -3019,
4020 => -2954,
4021 => -2888,
4022 => -2823,
4023 => -2757,
4024 => -2692,
4025 => -2626,
4026 => -2561,
4027 => -2495,
4028 => -2429,
4029 => -2364,
4030 => -2298,
4031 => -2233,
4032 => -2167,
4033 => -2101,
4034 => -2036,
4035 => -1970,
4036 => -1904,
4037 => -1839,
4038 => -1773,
4039 => -1707,
4040 => -1642,
4041 => -1576,
4042 => -1510,
4043 => -1444,
4044 => -1379,
4045 => -1313,
4046 => -1247,
4047 => -1181,
4048 => -1116,
4049 => -1050,
4050 => -984,
4051 => -918,
4052 => -852,
4053 => -787,
4054 => -721,
4055 => -655,
4056 => -589,
4057 => -523,
4058 => -457,
4059 => -392,
4060 => -326,
4061 => -260,
4062 => -194,
4063 => -128,
4064 => -62,
4065 => 4,
4066 => 69,
4067 => 135,
4068 => 201,
4069 => 267,
4070 => 333,
4071 => 399,
4072 => 465,
4073 => 531,
4074 => 597,
4075 => 663,
4076 => 729,
4077 => 794,
4078 => 860,
4079 => 926,
4080 => 992,
4081 => 1058,
4082 => 1124,
4083 => 1190,
4084 => 1256,
4085 => 1322,
4086 => 1388,
4087 => 1454,
4088 => 1520,
4089 => 1586,
4090 => 1652,
4091 => 1718,
4092 => 1784,
4093 => 1850,
4094 => 1916,
4095 => 1982
);


	COMPONENT spi_master is
			PORT (
	      clk_in : in  STD_LOGIC; --
			Data1 : in  std_logic_vector(11 DOWNTO 0);
			Data2 : in  STD_LOGIC_VECTOR(11 DOWNTO 0);
			
			CS_spi : out std_logic;
			CLK_spi : out std_logic;
			MOSI1_spi  : out std_logic;
			MOSI2_spi  : out std_logic
	  );
	END COMPONENT;	
	
	COMPONENT filter is
		PORT (
		clk : in  STD_LOGIC; --
		clk_enable : in  std_logic;
		reset : in  STD_LOGIC;
		
		filter_in : in std_logic_vector(11 downto 0);
		filter_out : out std_logic_vector(11 downto 0)
	  );
	END COMPONENT;	
	
	COMPONENT ADC_priem is
			PORT (
	      clk_in : in  STD_LOGIC; 
			
			CS_spi : out std_logic;
			CLK_spi : out std_logic;
			MOSI1_spi  : in std_logic;
			MOSI2_spi  : in std_logic;
			
			DataADC : out std_logic_vector(11 downto 0)
	  );
	END COMPONENT;	

begin
	
	led <= "10101010";
	
	process(clk_da2)
	begin
		if (clk_da2'event and clk_da2 = '1') then
			if (i = 4095) then
				i<=0;
			else i <= i + 1;	
			end if;
		end if;	
	end process;

--	process(clk_da2)
--	begin
--		if (clk_da2'event and clk_da2 = '1') then
--			ink <= 1;
--			if (pila + ink > 4095) then
--				pila <= 0;
--			else pila <= pila + ink;
--			end if;
--		end if;
--	end process;	
	
	Data1 <= std_logic_vector(to_unsigned(sin_array(i),12));
	Data2 <= std_logic_vector(to_unsigned(sin_array(i),12));
	
	process(clk)
	begin
	if (clk'event and clk = '1') then
		if (switch(0) = '1') then 
			RES_out <= ADC1; 
		else RES_out <= ADC; 
		end if;
	end if;	
	end process;
	
	spi : spi_master
		port map(
            clk_in => clk, -- ~5.3 Hz
				Data1 =>  Res_out,
				Data2 => Data2,			
				
				CS_spi => nSync,
				CLK_spi => CLK_DAC,
				MOSI1_spi => D1,
				MOSI2_spi => D2
		);
	
--	cs_sp <= cs_spi;

	ADCrwfgwg : ADC_priem
		port map(
            clk_in => clk, -- 		
				
				CS_spi => nSync_ADC,
				CLK_spi => CLK_ADC,
				MOSI1_spi => DataADC,--D2
				MOSI2_spi => DataADC2,
				
				DataADC => ADC
		);
		
	filtr_kih : filter
		port map(
		clk => clk_da2,
		clk_enable => switch(1),
		reset => switch(2),
		filter_in => ADC,
		filter_out => ADC1
		);
	
	process (clk)
	--suda cnt
	begin
		if rising_edge(clk) then	
			if cnt = 1151 then 
				cnt <= 0;
				clk_da2 <= not clk_da2;
			else 
				cnt <= cnt + 1;
			end if;
		end if;
	end process;	

end Behavioral;

